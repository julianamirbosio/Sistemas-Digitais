use ieee.std_logic_1164.all;

entity fibonacci is
    generic(width: positive := 16);
    port(
		-- control inputs
        clock, clear: in std_logic;
		iniciar: in std_logic;
		-- control outputs
		pronto: out std_logic;
		-- data inputs
        n: in std_logic_vector(width-1 downto 0);
		-- data outputs
        nterm: out std_logic_vector(width-1 downto 0)
    );
end entity;

architecture structure of fibonacci is
    component fibonacciControlBlock is
        port(
            clock, clear: in std_logic;
            ctrl1, ctrl2, ctrl3, ctrl4, ctrl5, ctrl6, ctrl7, ctrl8, ctrl9: out std_logic;
            stt1, stt2: in std_logic;
			iniciar: in std_logic;
			pronto: out std_logic
        );
    end component;
    
    component fibonacciOperatingBlock is
        generic(width: positive);
        port(
            clock, clear: in std_logic;
            ctrl1, ctrl2, ctrl3, ctrl4, ctrl5, ctrl6, ctrl7, ctrl8, ctrl9: in std_logic;
            stt1, stt2: out std_logic;
            n: in std_logic_vector(width-1 downto 0);
            nterm: out std_logic_vector(width-1 downto 0)
        );
    end component;

    signal  -- COMPLETE
begin
    BC: fibonacciControlBlock port map(--COMPLETE);
    BO: fibonacciOperatingBlock generic map(width) port map(--COMPLETE);
end architecture;
